module sine_float(theta,sign,exponenet,theta_out);

input [31:0] theta;
real pi_mantissa 1.5707963267948966
real two_pi_exponent 2

endmodule